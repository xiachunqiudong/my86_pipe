`include "define.v"

module execute_reg();


endmodule